library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity gen_mux is
	generic (BREITE : positive := 8);
end entity gen_mux;

architecture RTL of gen_mux is
	
begin

end architecture RTL;
